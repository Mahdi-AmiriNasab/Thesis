** Profile: "SCHEMATIC1-switch_sim"  [ D:\Thesis\pspice\test-SCHEMATIC1-switch_sim.sim ] 

** Creating circuit file "test-SCHEMATIC1-switch_sim.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1 0 1e-3 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\test-SCHEMATIC1.net" 


.END
